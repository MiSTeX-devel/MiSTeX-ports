-- megafunction wizard: %RAM: 2-PORT%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: altdpram 

-- ============================================================
-- File Name: cx4cache.vhd
-- Megafunction Name(s):
-- 			altdpram
--
-- Simulation Library Files(s):
-- 			altera_mf
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 13.1.4 Build 182 03/12/2014 SJ Full Version
-- ************************************************************


--Copyright (C) 1991-2014 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;


ENTITY cx4cache IS
	PORT
	(
		clock		: IN STD_LOGIC ;
		data		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		rdaddress	: IN STD_LOGIC_VECTOR (8 DOWNTO 0);
		wraddress	: IN STD_LOGIC_VECTOR (8 DOWNTO 0);
		wren		: IN STD_LOGIC  := '0';
		q		    : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
	);
END cx4cache;


ARCHITECTURE SYN OF cx4cache IS
constant addr_width : positive := 9;
constant data_width : positive := 8;

constant DEPTH        :  positive := 2**addr_width;
subtype  word_t	      is std_logic_vector(data_width - 1 downto 0);
type	 ram_t		  is array(0 to DEPTH - 1) of word_t;
signal   ram          :  ram_t;

begin
process (clock)
begin
	if rising_edge(clock) then
		if wren = '1' then
			ram(to_integer(unsigned(wraddress))) <= data;
		end if;
		q <= ram(to_integer(unsigned(rdaddress)));
	end if;
end process;

END SYN;
